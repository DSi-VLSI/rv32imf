// Module to perform a fancy shift and find the first '1' from the left
module pa_fdsu_ff1 (
    fanc_shift_num,  // Output: Shifted fraction number
    frac_bin_val,  // Output: Binary value indicating position of first '1'
    frac_num  // Input: 52-bit fraction number
);

  input [51:0] frac_num;  // Input: 52-bit fraction number
  output [51:0] fanc_shift_num;  // Output: Shifted fraction number
  output [12:0] frac_bin_val;  // Output: Binary value for first '1' position

  reg  [51:0] fanc_shift_num;  // Register for shifted fraction number
  reg  [12:0] frac_bin_val;  // Register for binary value of first '1'

  wire [51:0] frac_num;  // Wire for input fraction number

  // Find the position of the first '1' from the left in frac_num
  always @(frac_num[51:0]) begin
    casez (frac_num[51:0])
      // If the first bit is '1'
      52'b1???????????????????????????????????????????????????: frac_bin_val[12:0] = 13'h0;
      // If the second bit is '1'
      52'b01??????????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1fff;
      // If the third bit is '1'
      52'b001?????????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ffe;
      // If the fourth bit is '1'
      52'b0001????????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ffd;
      // If the fifth bit is '1'
      52'b00001???????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ffc;
      // If the sixth bit is '1'
      52'b000001??????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ffb;
      // If the seventh bit is '1'
      52'b0000001?????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ffa;
      // If the eighth bit is '1'
      52'b00000001????????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff9;
      // If the ninth bit is '1'
      52'b000000001???????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff8;
      // If the tenth bit is '1'
      52'b0000000001??????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff7;
      // If the eleventh bit is '1'
      52'b00000000001?????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff6;
      // If the twelfth bit is '1'
      52'b000000000001????????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff5;
      // If the thirteenth bit is '1'
      52'b0000000000001???????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff4;
      // If the fourteenth bit is '1'
      52'b00000000000001??????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff3;
      // If the fifteenth bit is '1'
      52'b000000000000001?????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff2;
      // If the sixteenth bit is '1'
      52'b0000000000000001????????????????????????????????????: frac_bin_val[12:0] = 13'h1ff1;
      // If the seventeenth bit is '1'
      52'b00000000000000001???????????????????????????????????: frac_bin_val[12:0] = 13'h1ff0;
      // If the eighteenth bit is '1'
      52'b000000000000000001??????????????????????????????????: frac_bin_val[12:0] = 13'h1fef;
      // If the nineteenth bit is '1'
      52'b0000000000000000001?????????????????????????????????: frac_bin_val[12:0] = 13'h1fee;
      // If the twentieth bit is '1'
      52'b00000000000000000001????????????????????????????????: frac_bin_val[12:0] = 13'h1fed;
      // If the twenty-first bit is '1'
      52'b000000000000000000001???????????????????????????????: frac_bin_val[12:0] = 13'h1fec;
      // If the twenty-second bit is '1'
      52'b0000000000000000000001??????????????????????????????: frac_bin_val[12:0] = 13'h1feb;
      // If the twenty-third bit is '1'
      52'b00000000000000000000001?????????????????????????????: frac_bin_val[12:0] = 13'h1fea;
      // If the twenty-fourth bit is '1'
      52'b000000000000000000000001????????????????????????????: frac_bin_val[12:0] = 13'h1fe9;
      // If the twenty-fifth bit is '1'
      52'b0000000000000000000000001???????????????????????????: frac_bin_val[12:0] = 13'h1fe8;
      // If the twenty-sixth bit is '1'
      52'b00000000000000000000000001??????????????????????????: frac_bin_val[12:0] = 13'h1fe7;
      // If the twenty-seventh bit is '1'
      52'b000000000000000000000000001?????????????????????????: frac_bin_val[12:0] = 13'h1fe6;
      // If the twenty-eighth bit is '1'
      52'b0000000000000000000000000001????????????????????????: frac_bin_val[12:0] = 13'h1fe5;
      // If the twenty-ninth bit is '1'
      52'b00000000000000000000000000001???????????????????????: frac_bin_val[12:0] = 13'h1fe4;
      // If the thirtieth bit is '1'
      52'b000000000000000000000000000001??????????????????????: frac_bin_val[12:0] = 13'h1fe3;
      // If the thirty-first bit is '1'
      52'b0000000000000000000000000000001?????????????????????: frac_bin_val[12:0] = 13'h1fe2;
      // If the thirty-second bit is '1'
      52'b00000000000000000000000000000001????????????????????: frac_bin_val[12:0] = 13'h1fe1;
      // If the thirty-third bit is '1'
      52'b000000000000000000000000000000001???????????????????: frac_bin_val[12:0] = 13'h1fe0;
      // If the thirty-fourth bit is '1'
      52'b0000000000000000000000000000000001??????????????????: frac_bin_val[12:0] = 13'h1fdf;
      // If the thirty-fifth bit is '1'
      52'b00000000000000000000000000000000001?????????????????: frac_bin_val[12:0] = 13'h1fde;
      // If the thirty-sixth bit is '1'
      52'b000000000000000000000000000000000001????????????????: frac_bin_val[12:0] = 13'h1fdd;
      // If the thirty-seventh bit is '1'
      52'b0000000000000000000000000000000000001???????????????: frac_bin_val[12:0] = 13'h1fdc;
      // If the thirty-eighth bit is '1'
      52'b00000000000000000000000000000000000001??????????????: frac_bin_val[12:0] = 13'h1fdb;
      // If the thirty-ninth bit is '1'
      52'b000000000000000000000000000000000000001?????????????: frac_bin_val[12:0] = 13'h1fda;
      // If the fortieth bit is '1'
      52'b0000000000000000000000000000000000000001????????????: frac_bin_val[12:0] = 13'h1fd9;
      // If the forty-first bit is '1'
      52'b00000000000000000000000000000000000000001???????????: frac_bin_val[12:0] = 13'h1fd8;
      // If the forty-second bit is '1'
      52'b000000000000000000000000000000000000000001??????????: frac_bin_val[12:0] = 13'h1fd7;
      // If the forty-third bit is '1'
      52'b0000000000000000000000000000000000000000001?????????: frac_bin_val[12:0] = 13'h1fd6;
      // If the forty-fourth bit is '1'
      52'b00000000000000000000000000000000000000000001????????: frac_bin_val[12:0] = 13'h1fd5;
      // If the forty-fifth bit is '1'
      52'b000000000000000000000000000000000000000000001???????: frac_bin_val[12:0] = 13'h1fd4;
      // If the forty-sixth bit is '1'
      52'b0000000000000000000000000000000000000000000001??????: frac_bin_val[12:0] = 13'h1fd3;
      // If the forty-seventh bit is '1'
      52'b00000000000000000000000000000000000000000000001?????: frac_bin_val[12:0] = 13'h1fd2;
      // If the forty-eighth bit is '1'
      52'b000000000000000000000000000000000000000000000001????: frac_bin_val[12:0] = 13'h1fd1;
      // If the forty-ninth bit is '1'
      52'b0000000000000000000000000000000000000000000000001???: frac_bin_val[12:0] = 13'h1fd0;
      // If the fiftieth bit is '1'
      52'b00000000000000000000000000000000000000000000000001??: frac_bin_val[12:0] = 13'h1fcf;
      // If the fifty-first bit is '1'
      52'b000000000000000000000000000000000000000000000000001?: frac_bin_val[12:0] = 13'h1fce;
      // If the fifty-second bit is '1'
      52'b0000000000000000000000000000000000000000000000000001: frac_bin_val[12:0] = 13'h1fcd;
      // If all bits are '0'
      52'b0000000000000000000000000000000000000000000000000000: frac_bin_val[12:0] = 13'h1fcc;
      // Default case
      default: frac_bin_val[12:0] = 13'h000;
    endcase
  end

  // Perform a fancy shift based on the position of the first '1'
  always @(frac_num[51:0]) begin
    casez (frac_num[51:0])
      // If the first bit is '1', no shift
      52'b1???????????????????????????????????????????????????:
      fanc_shift_num[51:0] = frac_num[51:0];
      // If the second bit is '1', shift left by 1
      52'b01??????????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[50:0], 1'b0};
      // If the third bit is '1', shift left by 2
      52'b001?????????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[49:0], 2'b0};
      // If the fourth bit is '1', shift left by 3
      52'b0001????????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[48:0], 3'b0};
      // If the fifth bit is '1', shift left by 4
      52'b00001???????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[47:0], 4'b0};
      // If the sixth bit is '1', shift left by 5
      52'b000001??????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[46:0], 5'b0};
      // If the seventh bit is '1', shift left by 6
      52'b0000001?????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[45:0], 6'b0};
      // If the eighth bit is '1', shift left by 7
      52'b00000001????????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[44:0], 7'b0};
      // If the ninth bit is '1', shift left by 8
      52'b000000001???????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[43:0], 8'b0};
      // If the tenth bit is '1', shift left by 9
      52'b0000000001??????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[42:0], 9'b0};
      // If the eleventh bit is '1', shift left by 10
      52'b00000000001?????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[41:0], 10'b0};
      // If the twelfth bit is '1', shift left by 11
      52'b000000000001????????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[40:0], 11'b0};
      // If the thirteenth bit is '1', shift left by 12
      52'b0000000000001???????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[39:0], 12'b0};
      // If the fourteenth bit is '1', shift left by 13
      52'b00000000000001??????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[38:0], 13'b0};
      // If the fifteenth bit is '1', shift left by 14
      52'b000000000000001?????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[37:0], 14'b0};
      // If the sixteenth bit is '1', shift left by 15
      52'b0000000000000001????????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[36:0], 15'b0};
      // If the seventeenth bit is '1', shift left by 16
      52'b00000000000000001???????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[35:0], 16'b0};
      // If the eighteenth bit is '1', shift left by 17
      52'b000000000000000001??????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[34:0], 17'b0};
      // If the nineteenth bit is '1', shift left by 18
      52'b0000000000000000001?????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[33:0], 18'b0};
      // If the twentieth bit is '1', shift left by 19
      52'b00000000000000000001????????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[32:0], 19'b0};
      // If the twenty-first bit is '1', shift left by 20
      52'b000000000000000000001???????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[31:0], 20'b0};
      // If the twenty-second bit is '1', shift left by 21
      52'b0000000000000000000001??????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[30:0], 21'b0};
      // If the twenty-third bit is '1', shift left by 22
      52'b00000000000000000000001?????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[29:0], 22'b0};
      // If the twenty-fourth bit is '1', shift left by 23
      52'b000000000000000000000001????????????????????????????:
      fanc_shift_num[51:0] = {frac_num[28:0], 23'b0};
      // If the twenty-fifth bit is '1', shift left by 24
      52'b0000000000000000000000001???????????????????????????:
      fanc_shift_num[51:0] = {frac_num[27:0], 24'b0};
      // If the twenty-sixth bit is '1', shift left by 25
      52'b00000000000000000000000001??????????????????????????:
      fanc_shift_num[51:0] = {frac_num[26:0], 25'b0};
      // If the twenty-seventh bit is '1', shift left by 26
      52'b000000000000000000000000001?????????????????????????:
      fanc_shift_num[51:0] = {frac_num[25:0], 26'b0};
      // If the twenty-eighth bit is '1', shift left by 27
      52'b0000000000000000000000000001????????????????????????:
      fanc_shift_num[51:0] = {frac_num[24:0], 27'b0};
      // If the twenty-ninth bit is '1', shift left by 28
      52'b00000000000000000000000000001???????????????????????:
      fanc_shift_num[51:0] = {frac_num[23:0], 28'b0};
      // If the thirtieth bit is '1', shift left by 29
      52'b000000000000000000000000000001??????????????????????:
      fanc_shift_num[51:0] = {frac_num[22:0], 29'b0};
      // If the thirty-first bit is '1', shift left by 30
      52'b0000000000000000000000000000001?????????????????????:
      fanc_shift_num[51:0] = {frac_num[21:0], 30'b0};
      // If the thirty-second bit is '1', shift left by 31
      52'b00000000000000000000000000000001????????????????????:
      fanc_shift_num[51:0] = {frac_num[20:0], 31'b0};
      // If the thirty-third bit is '1', shift left by 32
      52'b000000000000000000000000000000001???????????????????:
      fanc_shift_num[51:0] = {frac_num[19:0], 32'b0};
      // If the thirty-fourth bit is '1', shift left by 33
      52'b0000000000000000000000000000000001??????????????????:
      fanc_shift_num[51:0] = {frac_num[18:0], 33'b0};
      // If the thirty-fifth bit is '1', shift left by 34
      52'b00000000000000000000000000000000001?????????????????:
      fanc_shift_num[51:0] = {frac_num[17:0], 34'b0};
      // If the thirty-sixth bit is '1', shift left by 35
      52'b000000000000000000000000000000000001????????????????:
      fanc_shift_num[51:0] = {frac_num[16:0], 35'b0};
      // If the thirty-seventh bit is '1', shift left by 36
      52'b0000000000000000000000000000000000001???????????????:
      fanc_shift_num[51:0] = {frac_num[15:0], 36'b0};
      // If the thirty-eighth bit is '1', shift left by 37
      52'b00000000000000000000000000000000000001??????????????:
      fanc_shift_num[51:0] = {frac_num[14:0], 37'b0};
      // If the thirty-ninth bit is '1', shift left by 38
      52'b000000000000000000000000000000000000001?????????????:
      fanc_shift_num[51:0] = {frac_num[13:0], 38'b0};
      // If the fortieth bit is '1', shift left by 39
      52'b0000000000000000000000000000000000000001????????????:
      fanc_shift_num[51:0] = {frac_num[12:0], 39'b0};
      // If the forty-first bit is '1', shift left by 40
      52'b00000000000000000000000000000000000000001???????????:
      fanc_shift_num[51:0] = {frac_num[11:0], 40'b0};
      // If the forty-second bit is '1', shift left by 41
      52'b000000000000000000000000000000000000000001??????????:
      fanc_shift_num[51:0] = {frac_num[10:0], 41'b0};
      // If the forty-third bit is '1', shift left by 42
      52'b0000000000000000000000000000000000000000001?????????:
      fanc_shift_num[51:0] = {frac_num[9:0], 42'b0};
      // If the forty-fourth bit is '1', shift left by 43
      52'b00000000000000000000000000000000000000000001????????:
      fanc_shift_num[51:0] = {frac_num[8:0], 43'b0};
      // If the forty-fifth bit is '1', shift left by 44
      52'b000000000000000000000000000000000000000000001???????:
      fanc_shift_num[51:0] = {frac_num[7:0], 44'b0};
      // If the forty-sixth bit is '1', shift left by 45
      52'b0000000000000000000000000000000000000000000001??????:
      fanc_shift_num[51:0] = {frac_num[6:0], 45'b0};
      // If the forty-seventh bit is '1', shift left by 46
      52'b00000000000000000000000000000000000000000000001?????:
      fanc_shift_num[51:0] = {frac_num[5:0], 46'b0};
      // If the forty-eighth bit is '1', shift left by 47
      52'b000000000000000000000000000000000000000000000001????:
      fanc_shift_num[51:0] = {frac_num[4:0], 47'b0};
      // If the forty-ninth bit is '1', shift left by 48
      52'b0000000000000000000000000000000000000000000000001???:
      fanc_shift_num[51:0] = {frac_num[3:0], 48'b0};
      // If the fiftieth bit is '1', shift left by 49
      52'b00000000000000000000000000000000000000000000000001??:
      fanc_shift_num[51:0] = {frac_num[2:0], 49'b0};
      // If the fifty-first bit is '1', shift left by 50
      52'b000000000000000000000000000000000000000000000000001?:
      fanc_shift_num[51:0] = {frac_num[1:0], 50'b0};
      // If the fifty-second bit is '1', shift left by 51
      52'b0000000000000000000000000000000000000000000000000001:
      fanc_shift_num[51:0] = {frac_num[0:0], 51'b0};
      // If all bits are '0', output all zeros
      52'b0000000000000000000000000000000000000000000000000000: fanc_shift_num[51:0] = {52'b0};
      // Default case
      default: fanc_shift_num[51:0] = {52'b0};
    endcase
  end

endmodule
