package rv32imf_apu_core_pkg;

  parameter int APU_NARGS_CPU = 3;
  parameter int APU_WOP_CPU = 6;
  parameter int APU_NDSFLAGS_CPU = 15;
  parameter int APU_NUSFLAGS_CPU = 5;

endpackage
